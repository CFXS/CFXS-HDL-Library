library ieee;
use ieee.std_logic_1164.all;

package Types is
end package;
